library ieee;
use ieee.std_logic_1164.all;

use work.config_pkg.all;

entity user_app is
    port (
        clk : in std_logic;
        rst : in std_logic;

        -- memory-map interface
        mmap_wr_en   : in  std_logic;
        mmap_wr_addr : in  std_logic_vector(MMAP_ADDR_RANGE);
        mmap_wr_data : in  std_logic_vector(MMAP_DATA_RANGE);
        mmap_rd_en   : in  std_logic;
        mmap_rd_addr : in  std_logic_vector(MMAP_ADDR_RANGE);
        mmap_rd_data : out std_logic_vector(MMAP_DATA_RANGE)
        );
end user_app;

architecture default of user_app is

  signal n      : std_logic_vector(31 downto 0);
  signal result : std_logic_vector(31 downto 0);
  signal done   : std_logic;
  signal go : std_logic;
begin
  
	-- connect memory map and fib entity
  mem_map : entity work.memory_map
    port map(
      clk     => clk,
      rst     => rst,
      wr_en   => mmap_wr_en,
      wr_addr => mmap_wr_addr,
      wr_data => mmap_wr_data,
      rd_en   => mmap_rd_en,
      rd_addr => mmap_rd_addr,
      rd_data => mmap_rd_data,
      go      => go,
      n       => n,
      result  => result,
      done    => done
    );
    
  fib : entity work.fib_fsmd
    generic map(
      width => 32
    )
    port map(
      clk => clk,
      rst => rst,
      go => go,
      n => n,
      done => done,
      result => result
    );

end default;
